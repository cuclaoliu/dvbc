//////////////////////////////////////////////////////////////////////////////
//
//	filename rsencoder.sv
//
//  The RS(204, 188)encode design file for DVB System. It includes two mode 
//		input iData stream frame structer. One is 188 bytes iData per frame with
//		1 synchronous byte, and the other is 204 bytes iData per frame with 1
//		synchronous byte and 16 bytes zero. The 16 bytes zero is added to the 
//		188 bytes iData before rs encode. The output iData stream will be 204 bytes
//		per frame. The first byte is the Synchronous byte. And the following 188
//		is the source iData to be transport. And the last 16 bytes are the error
//		correct code for the 188 bytes witch is generated by this module and added
//		or filled to the tail of the input iData stream.
//
//////////////////////////////////////////////////////////////////////-
//	rev: 2.0
//	author: Liuchy
//	date: May 9, 2008
////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ns

module rsenc(
	iClk,
	iClrn,
	iData,
	iValid,
	iPSync,
	iCheck,
	oData,
	oPSync, 
	oValid
	);
	
	output logic[7:0] oData = 8'b0;
	output logic oPSync = 1'b0;
	output logic oValid = 1'b0;
	input iClk, iClrn, iCheck;
	input iPSync, iValid;
	input[7:0] iData;
	
	//	Declare the registers
	logic[7:0] data_reg [15:0];
	logic IsParity;
	logic[7:0] multiplier;
	logic[7:0] multiplier_alpha;
	logic[7:0] product[15:0];
	logic[7:0] product_x[15:0];
	byte unsigned bytescnt;
	
	assign multiplier = iCheck?8'b0:(iData^data_reg[15]);
	integer loop_v;//for for statement
	
	always_ff @(posedge iClk or negedge iClrn) begin
		if(!iClrn) begin
			for (loop_v=0; loop_v<=15; loop_v=loop_v+1) begin
				data_reg[loop_v] <= #1 8'b0;
			end
		end
		else if(iValid) begin
			data_reg[0] <= #1 product_x[0];
			for (loop_v=1; loop_v<=15; loop_v=loop_v+1) begin
				//if(iPSync)
				//	data_reg[loop_v] <= #1 8'd0;
				//else
					data_reg[loop_v] <= #1 data_reg[loop_v-1] ^ product_x[loop_v];
			end
			if (iCheck)
				oData <= #1 data_reg[15];
			else
				oData <= #1 iData;
		end
	end
	
	always_ff @(posedge iClk or negedge iClrn) begin
		if (!iClrn) begin
			oValid <= #1 1'b0;
			oPSync <= #1 1'b0;
			bytescnt <= #1 8'd0;
			//IsParity <= #1 1'b0;
		end
		else begin
			oValid <= #1 iValid;
			oPSync <= #1 iPSync;
			if(iPSync & iValid) begin
				bytescnt <= #1 8'd1;
				//IsParity <= #1 1'b0;
			end
			else if(iValid) begin
				if(bytescnt < 203)
					bytescnt <= #1 bytescnt + 8'd1;
				else
					bytescnt <= #1 8'd0;
			end
		end
	end
	
	canonical2dual canonical2dual_inst(
		.canonical(multiplier), .dual(multiplier_alpha));
		
	//	Declare the lookup table for a(n)*g(r)
	//	The coefficient of generator polynomial is 
	//		g[15..0] : 59,13,104,189,68,209,30,8,163,65,41,229,98,50,36,59
	//		g[15]=g[0]=59 will share just one lut result.
	multiplier_120 multiplier00(
		.in(multiplier_alpha), .out(product[0]));
	dual2canonical dual2canonical00(
		.dual(product[0]), .canonical(product_x[0]));
	multiplier_225 multiplier01(
		.in(multiplier_alpha), .out(product[1]));
	dual2canonical dual2canonical01(
		.dual(product[1]), .canonical(product_x[1]));
	multiplier_194 multiplier02(
		.in(multiplier_alpha), .out(product[2]));
	dual2canonical dual2canonical02(
		.dual(product[2]), .canonical(product_x[2]));
	multiplier_182 multiplier03(
		.in(multiplier_alpha), .out(product[3]));
	dual2canonical dual2canonical03(
		.dual(product[3]), .canonical(product_x[3]));
	multiplier_169 multiplier04(
		.in(multiplier_alpha), .out(product[4]));
	dual2canonical dual2canonical04(
		.dual(product[4]), .canonical(product_x[4]));
	multiplier_147 multiplier05(
		.in(multiplier_alpha), .out(product[5]));
	dual2canonical dual2canonical05(
		.dual(product[5]), .canonical(product_x[5]));
	multiplier_191 multiplier06(
		.in(multiplier_alpha), .out(product[6]));
	dual2canonical dual2canonical06(
		.dual(product[6]), .canonical(product_x[6]));
	multiplier_91 multiplier07(
		.in(multiplier_alpha), .out(product[7]));
	dual2canonical dual2canonical07(
		.dual(product[7]), .canonical(product_x[7]));
	multiplier_3 multiplier08(
		.in(multiplier_alpha), .out(product[8]));
	dual2canonical dual2canonical08(
		.dual(product[8]), .canonical(product_x[8]));
	multiplier_76 multiplier09(
		.in(multiplier_alpha), .out(product[9]));
	dual2canonical dual2canonical09(
		.dual(product[9]), .canonical(product_x[9]));
	multiplier_161 multiplier10(
		.in(multiplier_alpha), .out(product[10]));
	dual2canonical dual2canonical10(
		.dual(product[10]), .canonical(product_x[10]));
	multiplier_102 multiplier11(
		.in(multiplier_alpha), .out(product[11]));
	dual2canonical dual2canonical11(
		.dual(product[11]), .canonical(product_x[11]));
	multiplier_109 multiplier12(
		.in(multiplier_alpha), .out(product[12]));
	dual2canonical dual2canonical12(
		.dual(product[12]), .canonical(product_x[12]));
	multiplier_107 multiplier13(
		.in(multiplier_alpha), .out(product[13]));
	dual2canonical dual2canonical13(
		.dual(product[13]), .canonical(product_x[13]));
	multiplier_104 multiplier14(
		.in(multiplier_alpha), .out(product[14]));
	dual2canonical dual2canonical14(
		.dual(product[14]), .canonical(product_x[14]));
	multiplier_120 multiplier15(
		.in(multiplier_alpha), .out(product[15]));
	dual2canonical dual2canonical15(
		.dual(product[15]), .canonical(product_x[15]));

endmodule

//////////////////////////////////////////////////////////////////////-
//	module name: canonical2dual
//
//	convert canonical basis to dual basis
//		w_tau0 = w_alpha7
//		w_tau1 = w_alpha6
//		w_tau2 = w_alpha5
//		w_tau3 = w_alpha4
//		w_tau4 = w_alpha7 + w_alpha3
//		w_tau5 = w_alpha7 + w_alpha6 + w_alpha2
//		w_tau6 = w_alpha7 + w_alpha6 + w_alpha5 + w_alpha1
//		w_tau7 = w_alpha6 + w_alpha5 + w_alpha4 + w_alpha0
//	note: the module-2 adder is implemented by ^.

module canonical2dual
(
	input[7:0] canonical,
	output[7:0] dual
);
	assign dual[0] = canonical[7];
	assign dual[1] = canonical[6];
	assign dual[2] = canonical[5];
	assign dual[3] = canonical[4];
	assign dual[4] = canonical[7] ^ canonical[3];
	assign dual[5] = canonical[7] ^ canonical[6] ^ canonical[2];
	assign dual[6] = canonical[7] ^ canonical[6] ^ canonical[5] ^ canonical[1];
	assign dual[7] = canonical[6] ^ canonical[5] ^ canonical[4] ^ canonical[0];
endmodule

//////////////////////////////////////////////////////////////////////-
//	module name: dual2canonical
//
//	convert dual basis to canonical basis
//		w_alpha7 = w_tau0
//		w_alpha6 = w_tau1
//		w_alpha5 = w_tau2
//		w_alpha4 = w_tau3
//		w_alpha3 = w_tau0 + w_tau4
//		w_alpha2 = w_tau0 + w_tau1 + w_tau5
//		w_alpha1 = w_tau0 + w_tau1 + w_tau2 + w_tau6
//		w_alpha0 = w_tau1 + w_tau2 + w_tau3 + w_tau7
//	note: the module-2 adder is implemented by ^.

module dual2canonical
(
	input [7:0]	dual,
	output[7:0] canonical
);

	assign canonical[0] = dual[1] ^ dual[2] ^ dual[3] ^ dual[7];
	assign canonical[1] = dual[0] ^ dual[1] ^ dual[2] ^ dual[6];
	assign canonical[2] = dual[0] ^ dual[1] ^ dual[5];
	assign canonical[3] = dual[0] ^ dual[4];
	assign canonical[4] = dual[3];
	assign canonical[5] = dual[2];
	assign canonical[6] = dual[1];
	assign canonical[7] = dual[0];
endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_120
//
//		w = uv
//		w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^120.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			w_tau0		0		0		1		1		1		0		1		1
//			w_tau1		0		1		1		1		0		1		1		0
//			w_tau2		1		1		1		0		1		1		0		0
//			w_tau3		1		1		0		0		0		1		0		1
//			w_tau4		1		0		0		1		0		1		1		1
//			w_tau5		0		0		1		1		0		0		1		1
//			w_tau6		0		1		1		0		0		1		1		0
//			w_tau7		1		1		0		0		1		1		0		0

module multiplier_120
(
	input[7:0] in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[1] = u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[2] ^ u_tau[1];
	assign w_tau[2] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[3] ^ u_tau[2];
	assign w_tau[3] = u_tau[7] ^ u_tau[6] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[4] = u_tau[7] ^ u_tau[4] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[5] = u_tau[5] ^ u_tau[4] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[6] = u_tau[6] ^ u_tau[5] ^ u_tau[2] ^ u_tau[1];
	assign w_tau[7] = u_tau[7] ^ u_tau[6] ^ u_tau[3] ^ u_tau[2];
	assign out = w_tau;

endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_225
//
//		w = uv
//		 w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^225.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			w_tau0		0		0		1		0		0		1		0		0
//			w_tau1		0		1		0		0		1		0		0		0
//			w_tau2		1		0		0		1		0		0		0		0
//			w_tau3		0		0		1		1		1		1		0		1
//			w_tau4		0		1		1		1		1		0		1		0
//			w_tau5		1		1		1		1		0		1		0		0
//			w_tau6		1		1		1		1		0		1		0		1
//			w_tau7		1		1		1		1		0		1		1		1

module multiplier_225
(
	input[7:0] in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[5] ^ u_tau[2];
	assign w_tau[1] = u_tau[6] ^ u_tau[3];
	assign w_tau[2] = u_tau[7] ^ u_tau[4];
	assign w_tau[3] = u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[4] = u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[1];
	assign w_tau[5] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[2];
	assign w_tau[6] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[7] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign out = w_tau;

endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_194
//
//		w = uv
//		w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^194.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			w_tau0		0		0		1		1		0		0		1		0
//			w_tau1		0		1		1		0		0		1		0		0
//			w_tau2		1		1		0		0		1		0		0		0
//			w_tau3		1		0		0		0		1		1		0		1
//			w_tau4		0		0		0		0		0		1		1		1
//			w_tau5		0		0		0		0		1		1		1		0
//			w_tau6		0		0		0		1		1		1		0		0
//			w_tau7		0		0		1		1		1		0		0		0

module multiplier_194
(
	input[7:0] in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[5] ^ u_tau[4] ^ u_tau[1];
	assign w_tau[1] = u_tau[6] ^ u_tau[5] ^ u_tau[2];
	assign w_tau[2] = u_tau[7] ^ u_tau[6] ^ u_tau[3];
	assign w_tau[3] = u_tau[7] ^ u_tau[3] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[4] = u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[5] = u_tau[3] ^ u_tau[2] ^ u_tau[1];
	assign w_tau[6] = u_tau[4] ^ u_tau[3] ^ u_tau[2];
	assign w_tau[7] = u_tau[5] ^ u_tau[4] ^ u_tau[3];
	assign out = w_tau[7:0];

endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_182
//
//		w = uv
//	a few steps
//		1. w_tau = u_tau * v; the logic convertion is base on a matlab program.
//		2. convert w_tau on dual basis to u on canonical basis.
//	for the multiplicator v = alpha^182.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			w_tau0		0		1		1		0		0		0		1		0
//			w_tau1		1		1		0		0		0		1		0		0
//			w_tau2		1		0		0		1		0		1		0		1
//			w_tau3		0		0		1		1		0		1		1		1
//			w_tau4		0		1		1		0		1		1		1		0
//			w_tau5		1		1		0		1		1		1		0		0
//			w_tau6		1		0		1		0		0		1		0		1
//			w_tau7		0		1		0		1		0		1		1		1

module multiplier_182
(
	input[7:0]	in,
	output[7:0] out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[6] ^ u_tau[5] ^ u_tau[1];
	assign w_tau[1] = u_tau[7] ^ u_tau[6] ^ u_tau[2];
	assign w_tau[2] = u_tau[7] ^ u_tau[4] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[3] = u_tau[5] ^ u_tau[4] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[4] = u_tau[6] ^ u_tau[5] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1];
	assign w_tau[5] = u_tau[7] ^ u_tau[6] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2];
	assign w_tau[6] = u_tau[7] ^ u_tau[5] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[7] = u_tau[6] ^ u_tau[4] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign out = w_tau;
	
endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_169
//
//		w = uv
//		w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^169.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			assign w_tau0		1		1		1		0		0		1		0		1
//			assign w_tau1		1		1		0		1		0		1		1		1
//			assign w_tau2		1		0		1		1		0		0		1		1
//			assign w_tau3		0		1		1		1		1		0		1		1
//			assign w_tau4		1		1		1		1		0		1		1		0
//			assign w_tau5		1		1		1		1		0		0		0		1
//			assign w_tau6		1		1		1		1		1		1		1		1
//			assign w_tau7		1		1		1		0		0		0		1		1

module multiplier_169
(
	input[7:0]	in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[1] = u_tau[7] ^ u_tau[6] ^ u_tau[4] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[2] = u_tau[7] ^ u_tau[5] ^ u_tau[4] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[3] = u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[4] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[2] ^ u_tau[1];
	assign w_tau[5] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[0];
	assign w_tau[6] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[7] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[1] ^ u_tau[0];
	assign out[7:0] = w_tau[7:0];

endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_147
//
//		w = uv
//		w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^147.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			assign w_tau0		0		0		1		0		1		0		0		1
//			assign w_tau1		0		1		0		1		0		0		1		0
//			assign w_tau2		1		0		1		0		0		1		0		0
//			assign w_tau3		0		1		0		1		0		1		0		1
//			assign w_tau4		1		0		1		0		1		0		1		0
//			assign w_tau5		0		1		0		0		1		0		0		1
//			assign w_tau6		1		0		0		1		0		0		1		0
//			assign w_tau7		0		0		1		1		1		0		0		1
module multiplier_147
(
	input[7:0]	in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[5] ^ u_tau[3] ^ u_tau[0];
	assign w_tau[1] = u_tau[6] ^ u_tau[4] ^ u_tau[1];
	assign w_tau[2] = u_tau[7] ^ u_tau[5] ^ u_tau[2];
	assign w_tau[3] = u_tau[6] ^ u_tau[4] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[4] = u_tau[7] ^ u_tau[5] ^ u_tau[3] ^ u_tau[1];
	assign w_tau[5] = u_tau[6] ^ u_tau[3] ^ u_tau[0];
	assign w_tau[6] = u_tau[7] ^ u_tau[4] ^ u_tau[1];
	assign w_tau[7] = u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[0];
	assign out[7:0] = w_tau[7:0];

endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_191
//
//		w = uv
//		w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^191.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			w_tau0		0		1		0		0		0		0		0		1
//			w_tau1		1		0		0		0		0		0		1		0
//			w_tau2		0		0		0		1		1		0		0		1
//			w_tau3		0		0		1		1		0		0		1		0
//			w_tau4		0		1		1		0		0		1		0		0
//			w_tau5		1		1		0		0		1		0		0		0
//			w_tau6		1		0		0		0		1		1		0		1
//			w_tau7		0		0		0		0		0		1		1		1
module multiplier_191
(
	input[7:0]	in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[6] ^ u_tau[0];
	assign w_tau[1] = u_tau[7] ^ u_tau[1];
	assign w_tau[2] = u_tau[4] ^ u_tau[3] ^ u_tau[0];
	assign w_tau[3] = u_tau[5] ^ u_tau[4] ^ u_tau[1];
	assign w_tau[4] = u_tau[6] ^ u_tau[5] ^ u_tau[2];
	assign w_tau[5] = u_tau[7] ^ u_tau[6] ^ u_tau[3];
	assign w_tau[6] = u_tau[7] ^ u_tau[3] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[7] = u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign out[7:0] = w_tau[7:0];

endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_91
//
//		w = uv
//		w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^91.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			assign w_tau0		1		0		1		0		0		0		1		1
//			assign w_tau1		0		1		0		1		1		0		1		1
//			assign w_tau2		1		0		1		1		0		1		1		0
//			assign w_tau3		0		1		1		1		0		0		0		1
//			assign w_tau4		1		1		1		0		0		0		1		0
//			assign w_tau5		1		1		0		1		1		0		0		1
//			assign w_tau6		1		0		1		0		1		1		1		1
//			assign w_tau7		0		1		0		0		0		0		1		1
module multiplier_91
(
	input[7:0]	in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[7] ^ u_tau[5] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[1] = u_tau[6] ^ u_tau[4] ^ u_tau[3] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[2] = u_tau[7] ^ u_tau[5] ^ u_tau[4] ^ u_tau[2] ^ u_tau[1];
	assign w_tau[3] = u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[0];
	assign w_tau[4] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[1];
	assign w_tau[5] = u_tau[7] ^ u_tau[6] ^ u_tau[4] ^ u_tau[3] ^ u_tau[0];
	assign w_tau[6] = u_tau[7] ^ u_tau[5] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[7] = u_tau[6] ^ u_tau[1] ^ u_tau[0];
	assign out[7:0] = w_tau[7:0];

endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_3
//
//		w = uv
//		w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^3.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			assign w_tau0		0		0		0		0		1		0		0		0
//			assign w_tau1		0		0		0		1		0		0		0		0
//			assign w_tau2		0		0		1		0		0		0		0		0
//			assign w_tau3		0		1		0		0		0		0		0		0
//			assign w_tau4		1		0		0		0		0		0		0		0
//			assign w_tau5		0		0		0		1		1		1		0		1
//			assign w_tau6		0		0		1		1		1		0		1		0
//			assign w_tau7		0		1		1		1		0		1		0		0
module multiplier_3
(
	input[7:0]	in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[3];
	assign w_tau[1] = u_tau[4];
	assign w_tau[2] = u_tau[5];
	assign w_tau[3] = u_tau[6];
	assign w_tau[4] = u_tau[7];
	assign w_tau[5] = u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[6] = u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[1];
	assign w_tau[7] = u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[2];
	assign out[7:0] = w_tau[7:0];

endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_76
//
//		w = uv
//		w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^76.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			assign w_tau0		0		0		0		1		1		1		1		0
//			assign w_tau1		0		0		1		1		1		1		0		0
//			assign w_tau2		0		1		1		1		1		0		0		0
//			assign w_tau3		1		1		1		1		0		0		0		0
//			assign w_tau4		1		1		1		1		1		1		0		1
//			assign w_tau5		1		1		1		0		0		1		1		1
//			assign w_tau6		1		1		0		1		0		0		1		1
//			assign w_tau7		1		0		1		1		1		0		1		1
module multiplier_76
(
	input[7:0]	in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1];
	assign w_tau[1] = u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2];
	assign w_tau[2] = u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3];
	assign w_tau[3] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[4];
	assign w_tau[4] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[5] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[6] = u_tau[7] ^ u_tau[6] ^ u_tau[4] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[7] = u_tau[7] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[1] ^ u_tau[0];
	assign out[7:0] = w_tau[7:0];

endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_161
//
//		w = uv
//		w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^161.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			assign w_tau0		1		1		0		1		0		0		0		1
//			assign w_tau1		1		0		1		1		1		1		1		1
//			assign w_tau2		0		1		1		0		0		0		1		1
//			assign w_tau3		1		1		0		0		0		1		1		0
//			assign w_tau4		1		0		0		1		0		0		0		1
//			assign w_tau5		0		0		1		1		1		1		1		1
//			assign w_tau6		0		1		1		1		1		1		1		0
//			assign w_tau7		1		1		1		1		1		1		0		0
module multiplier_161
(
	input[7:0]	in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[7] ^ u_tau[6] ^ u_tau[4] ^ u_tau[0];
	assign w_tau[1] = u_tau[7] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[2] = u_tau[6] ^ u_tau[5] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[3] = u_tau[7] ^ u_tau[6] ^ u_tau[2] ^ u_tau[1];
	assign w_tau[4] = u_tau[7] ^ u_tau[4] ^ u_tau[0];
	assign w_tau[5] = u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[6] = u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1];
	assign w_tau[7] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2];
	assign out[7:0] = w_tau[7:0];

endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_102
//
//		w = uv
//		w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^102.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			assign w_tau0		0		1		0		0		0		1		0		0
//			assign w_tau1		1		0		0		0		1		0		0		0
//			assign w_tau2		0		0		0		0		1		1		0		1
//			assign w_tau3		0		0		0		1		1		0		1		0
//			assign w_tau4		0		0		1		1		0		1		0		0
//			assign w_tau5		0		1		1		0		1		0		0		0
//			assign w_tau6		1		1		0		1		0		0		0		0
//			assign w_tau7		1		0		1		1		1		1		0		1
module multiplier_102
(
	input[7:0]	in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[6] ^ u_tau[2];
	assign w_tau[1] = u_tau[7] ^ u_tau[3];
	assign w_tau[2] = u_tau[3] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[3] = u_tau[4] ^ u_tau[3] ^ u_tau[1];
	assign w_tau[4] = u_tau[5] ^ u_tau[4] ^ u_tau[2];
	assign w_tau[5] = u_tau[6] ^ u_tau[5] ^ u_tau[3];
	assign w_tau[6] = u_tau[7] ^ u_tau[6] ^ u_tau[4];
	assign w_tau[7] = u_tau[7] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[0];
	assign out[7:0] = w_tau[7:0];

endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_109
//
//		w = uv
//		w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^109.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			assign w_tau0		1		0		1		1		1		1		0		1
//			assign w_tau1		0		1		1		0		0		1		1		1
//			assign w_tau2		1		1		0		0		1		1		1		0
//			assign w_tau3		1		0		0		0		0		0		0		1
//			assign w_tau4		0		0		0		1		1		1		1		1
//			assign w_tau5		0		0		1		1		1		1		1		0
//			assign w_tau6		0		1		1		1		1		1		0		0
//			assign w_tau7		1		1		1		1		1		0		0		0
module multiplier_109
(
	input[7:0]	in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[7] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[1] = u_tau[6] ^ u_tau[5] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[2] = u_tau[7] ^ u_tau[6] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1];
	assign w_tau[3] = u_tau[7] ^ u_tau[0];
	assign w_tau[4] = u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[5] = u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1];
	assign w_tau[6] = u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2];
	assign w_tau[7] = u_tau[7] ^ u_tau[6] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3];
	assign out[7:0] = w_tau[7:0];

endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_107
//
//		w = uv
//		w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^107.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			assign w_tau0		0		1		1		0		1		0		0		0
//			assign w_tau1		1		1		0		1		0		0		0		0
//			assign w_tau2		1		0		1		1		1		1		0		1
//			assign w_tau3		0		1		1		0		0		1		1		1
//			assign w_tau4		1		1		0		0		1		1		1		0
//			assign w_tau5		1		0		0		0		0		0		0		1
//			assign w_tau6		0		0		0		1		1		1		1		1
//			assign w_tau7		0		0		1		1		1		1		1		0
module multiplier_107
(
	input[7:0]	in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[6] ^ u_tau[5] ^ u_tau[3];
	assign w_tau[1] = u_tau[7] ^ u_tau[6] ^ u_tau[4];
	assign w_tau[2] = u_tau[7] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[3] = u_tau[6] ^ u_tau[5] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[4] = u_tau[7] ^ u_tau[6] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1];
	assign w_tau[5] = u_tau[7] ^ u_tau[0];
	assign w_tau[6] = u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[7] = u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1];
	assign out[7:0] = w_tau[7:0];

endmodule

//////////////////////////////////////////////////////////////////////////////-
//
//	module name: multiplier_104
//
//		w = uv
//		w_tau = u_tau * v; the logic convertion is base on a matlab program.
//	for the multiplicator v = alpha^104.
//		+element	u_tau7	u_tau6	u_tau5	u_tau4	u_tau3	u_tau2	u_tau1	u_tau0
//			assign w_tau0		0		0		0		0		1		1		0		1
//			assign w_tau1		0		0		0		1		1		0		1		0
//			assign w_tau2		0		0		1		1		0		1		0		0
//			assign w_tau3		0		1		1		0		1		0		0		0
//			assign w_tau4		1		1		0		1		0		0		0		0
//			assign w_tau5		1		0		1		1		1		1		0		1
//			assign w_tau6		0		1		1		0		0		1		1		1
//			assign w_tau7		1		1		0		0		1		1		1		0
module multiplier_104
(
	input[7:0]	in,
	output[7:0]	out
);

	logic[7:0] u_tau;
	logic[7:0] w_tau;
	assign u_tau = in;
	assign w_tau[0] = u_tau[3] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[1] = u_tau[4] ^ u_tau[3] ^ u_tau[1];
	assign w_tau[2] = u_tau[5] ^ u_tau[4] ^ u_tau[2];
	assign w_tau[3] = u_tau[6] ^ u_tau[5] ^ u_tau[3];
	assign w_tau[4] = u_tau[7] ^ u_tau[6] ^ u_tau[4];
	assign w_tau[5] = u_tau[7] ^ u_tau[5] ^ u_tau[4] ^ u_tau[3] ^ u_tau[2] ^ u_tau[0];
	assign w_tau[6] = u_tau[6] ^ u_tau[5] ^ u_tau[2] ^ u_tau[1] ^ u_tau[0];
	assign w_tau[7] = u_tau[7] ^ u_tau[6] ^ u_tau[3] ^ u_tau[2] ^ u_tau[1];
	assign out[7:0] = w_tau[7:0];

endmodule